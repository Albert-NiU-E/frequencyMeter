LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY GATESIGNAL IS
PORT (
		LOCK    : OUT STD_LOGIC;
		GOUT    : OUT STD_LOGIC;
		CLEAR   : OUT STD_LOGIC;
		S1      : IN  STD_LOGIC;
		S2      : IN  STD_LOGIC;
		CLK     : IN  STD_LOGIC
		);
END GATESIGNAL;

ARCHITECTURE ARCHITECTURE_GATE OF GATESIGNAL IS

BEGIN
--======十分频计数========--
	PROCESS(CLK)
	VARIABLE COUNT:INTEGER:=0;
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			IF (S2 = '0' AND S1 = '0') THEN
				IF (COUNT > 10) THEN
					COUNT := 0;
				ELSE COUNT := COUNT + 1;
				END IF;
			END IF;
		END IF;
	END PROCESS;
--=====锁存信号========--
PROCESS(CLK)
VARIABLE COUNT:INTEGER:=0;
BEGIN
	IF(CLK'EVENT AND CLK = '1') THEN
		IF(COUNT=0) THEN
			LOCK <= '0';
		ELSE 
			LOCK <= '1';
		END IF;
	END IF;
END PROCESS;
--======清零信号========--
PROCESS(CLK)
VARIABLE COUNT:INTEGER:=0;
BEGIN
	IF (CLK'EVENT AND CLK = '1') THEN
		IF (COUNT >= 1) THEN
			CLEAR <= '0';
		ELSE
			CLEAR <= '1';
		END IF;
	END IF;
END PROCESS;

--=====GOUT作为使能端计数=======--
PROCESS(CLK)
VARIABLE COUNT:INTEGER:=0;
BEGIN
	IF (CLK'EVENT AND CLK = '1') THEN
		IF(COUNT >1) THEN
			GOUT <= '1';
		ELSE
			GOUT <= '0';
		END IF;
	END IF;
END PROCESS;

END ARCHITECTURE_GATE;