LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SECONDS IS
PORT (
		SECONDS    : OUT STD_LOGIC;
		CLK       : IN  STD_LOGIC
		); 
END SECONDS;

ARCHITECTURE ARCHITECTURE_SECONDS OF SECONDS IS
SIGNAL SEC: STD_LOGIC;
BEGIN
	PROCESS(CLK)--200Hz分频
	VARIABLE COUNT_SEC:INTEGER:=0;
	BEGIN
		IF(CLK'EVENT AND CLK = '1') THEN
			COUNT_SEC:=COUNT_SEC + 1;
			IF(COUNT_SEC<25000001) THEN 
				SEC <= '1';
			ELSIF(COUNT_SEC < 50000001) THEN 
				SEC <= '0';
			ELSE COUNT_SEC:=0;
			END IF;
		END IF;
		SECONDS<=SEC;
	END PROCESS;
END ARCHITECTURE_SECONDS;