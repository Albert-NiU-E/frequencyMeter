LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY LOCK IS
	PORT (
	LOCK    : IN STD_LOGIC;
	Q1      : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	Q2      : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	Q3      : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	QOUT    : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
	HZERO   : OUT STD_LOGIC:='0'
	);
END LOCK;

ARCHITECTURE ARCHITECTURE_LOCK OF LOCK IS
	SIGNAL Q321 : STD_LOGIC_VECTOR(11 DOWNTO 0);
BEGIN


--=======锁存========--
	PROCESS(LOCK)
	BEGIN
		IF(LOCK'EVENT AND LOCK = '0') THEN
			Q321 <= (Q3 & Q2 & Q1);
			QOUT <= Q321;
		END IF;
	END PROCESS;
	
	
--====判断是否有高位零，有就让HZERO使能传给AUTO===
	PROCESS(LOCK)
	BEGIN
		IF(LOCK'EVENT AND LOCK = '0') THEN
			IF(Q3 = "0000") THEN
				HZERO <= '1';
			ELSE
				HZERO <= '0';
			END IF;
		END IF;
	END PROCESS;
END ARCHITECTURE_LOCK;
		