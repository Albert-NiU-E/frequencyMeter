LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TESTIN IS
PORT(
	TEST  :   IN STD_LOGIC;
	S2    :   IN STD_LOGIC;
	CP    :   OUT STD_LOGIC
);
END TESTIN;

ARCHITECTURE ARCHITECTURE_TESTIN OF TESTIN IS
SIGNAL MODE : STD_LOGIC;
BEGIN
--=====高频十分频设计=========--
	PROCESS(TEST)
		VARIABLE COUNT_10H :INTEGER:= 0;
	BEGIN
			IF(TEST'EVENT AND TEST = '1') THEN
				COUNT_10H := COUNT_10H + 1;
				IF ( COUNT_10H <= 5 ) THEN 
					MODE <= '1';
				ELSIF (COUNT_10H <= 10) THEN
					MODE <= '0';
				ELSE COUNT_10H := 0;
				END IF;
			END IF;
	END PROCESS;

--=======模式选择==========--
PROCESS(TEST,S2)
BEGIN
	IF (S2 = '1') THEN
		CP <= MODE;
	ELSE
		CP <= TEST;
	END IF;
END PROCESS;

END ARCHITECTURE_TESTIN;